library verilog;
use verilog.vl_types.all;
entity MC68K is
    port(
        altera_reserved_tms: in     vl_logic;
        altera_reserved_tck: in     vl_logic;
        altera_reserved_tdi: in     vl_logic;
        altera_reserved_tdo: out    vl_logic;
        CPUClock        : out    vl_logic;
        CLK_50Mhz       : in     vl_logic;
        sdram_cke       : out    vl_logic;
        RESET_Key0_L    : in     vl_logic;
        AS_L            : out    vl_logic;
        UDS_L           : out    vl_logic;
        DataBusOut      : out    vl_logic_vector(15 downto 0);
        FlashData       : inout  vl_logic_vector(7 downto 0);
        LDS_L           : out    vl_logic;
        Bus_Request_SW8_H: in     vl_logic;
        DataBusIn       : out    vl_logic_vector(15 downto 0);
        SRam_Data       : inout  vl_logic_vector(15 downto 0);
        InPortA         : in     vl_logic_vector(7 downto 0);
        InPortB         : in     vl_logic_vector(7 downto 0);
        InPortC         : in     vl_logic_vector(7 downto 0);
        InPortE         : in     vl_logic_vector(7 downto 0);
        RS232_RxData    : in     vl_logic;
        Trace_Request_Key3_L: in     vl_logic;
        IRQ4_Key1_L     : in     vl_logic;
        IRQ2_Key2_L     : in     vl_logic;
        DMA_DataOut     : out    vl_logic_vector(15 downto 0);
        sdram_dq        : inout  vl_logic_vector(15 downto 0);
        sdram_cs_n      : out    vl_logic;
        sdram_ras_n     : out    vl_logic;
        sdram_cas_n     : out    vl_logic;
        sdram_we_n      : out    vl_logic;
        RomSelect_H     : out    vl_logic;
        Dtack_L         : out    vl_logic;
        sdram_clock     : out    vl_logic;
        LCD_RW          : out    vl_logic;
        CPU_RW          : out    vl_logic;
        LCD_E           : out    vl_logic;
        LCD_RS          : out    vl_logic;
        horiz_sync_out  : out    vl_logic;
        vert_sync_out   : out    vl_logic;
        SRam_OE_L       : out    vl_logic;
        SRam_CE_L       : out    vl_logic;
        SRam_WE_L       : out    vl_logic;
        SRam_LB_L       : out    vl_logic;
        SRam_UB_L       : out    vl_logic;
        ResetOut        : out    vl_logic;
        DramDtack_L     : out    vl_logic;
        FlashOE_L       : out    vl_logic;
        FlashWE_L       : out    vl_logic;
        FlashReset_L    : out    vl_logic;
        FlashCE_L       : out    vl_logic;
        DramSelect_H    : out    vl_logic;
        RS232_TxData    : out    vl_logic;
        OnChipRamSelect_H: out    vl_logic;
        BG_L            : out    vl_logic;
        LCD_Contrast_DE1: out    vl_logic;
        LCD_BLON_DE2    : out    vl_logic;
        LCD_ON_DE2      : out    vl_logic;
        UDS_OUT_L       : out    vl_logic;
        LDS_OUT_L       : out    vl_logic;
        RW_OUT          : out    vl_logic;
        AS_OUT_L        : out    vl_logic;
        BR_L            : out    vl_logic;
        BGACK_L         : out    vl_logic;
        VideoDac_Sync_L : out    vl_logic;
        VideoDac_Clock  : out    vl_logic;
        VideoDAC_Blank_L: out    vl_logic;
        SRamSelect_H    : out    vl_logic;
        Address_OUT     : out    vl_logic_vector(31 downto 0);
        AddressBus      : out    vl_logic_vector(31 downto 0);
        BlueOut         : out    vl_logic_vector(9 downto 0);
        FlashAddress    : out    vl_logic_vector(21 downto 0);
        GreenLEDS       : out    vl_logic_vector(7 downto 0);
        GreenOut        : out    vl_logic_vector(9 downto 0);
        HexDisplay0     : out    vl_logic_vector(6 downto 0);
        HexDisplay1     : out    vl_logic_vector(6 downto 0);
        HexDisplay2     : out    vl_logic_vector(6 downto 0);
        HexDisplay3     : out    vl_logic_vector(6 downto 0);
        HexDisplay4     : out    vl_logic_vector(6 downto 0);
        HexDisplay5     : out    vl_logic_vector(6 downto 0);
        HexDisplay6     : out    vl_logic_vector(6 downto 0);
        HexDisplay7     : out    vl_logic_vector(6 downto 0);
        LCDDataOut      : out    vl_logic_vector(7 downto 0);
        OutPortE        : out    vl_logic_vector(7 downto 0);
        RedLEDSA        : out    vl_logic_vector(7 downto 0);
        RedLEDSB        : out    vl_logic_vector(7 downto 0);
        RedLEDSC        : out    vl_logic_vector(7 downto 0);
        RedOut          : out    vl_logic_vector(9 downto 0);
        sdram_a         : out    vl_logic_vector(11 downto 0);
        sdram_ba        : out    vl_logic_vector(1 downto 0);
        sdram_dqm       : out    vl_logic_vector(1 downto 0);
        SRamAddress     : out    vl_logic_vector(17 downto 0)
    );
end MC68K;
