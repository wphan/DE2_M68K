LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all ;

-- 5 by 7 pixel ASCii character generator rom

entity CharacterGenRom5x7 is
	Port (
	
		Address	: in std_logic_Vector(9 downto 0);		-- 1024 locations 
		DataOut  : out std_logic_vector(7 downto 0)		-- a byte
	);
end ;


architecture bhvr of CharacterGenRom5x7 is
	type CharRom5x7 is array ( 0 to 1023) of std_logic_vector(7 downto 0);
	constant MyRom : CharRom5x7 := 
						(
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",	 		--  ' '
								X"00",X"04",X"04",X"04",X"04",X"00",X"00",X"04", 			--  '!'
								X"00",X"0a",X"0a",X"0a",X"00",X"00",X"00",X"00", 			--  '"'
								X"00",X"0a",X"0a",X"1f",X"0a",X"1f",X"0a",X"0a", 			--  '#'
								X"00",X"04",X"0f",X"14",X"0e",X"05",X"1e",X"04", 			--  '$'
								X"00",X"18",X"19",X"02",X"04",X"08",X"13",X"13", 			--  '%'
								X"00",X"0c",X"12",X"14",X"08",X"15",X"12",X"0d", 			--  '&'
								X"00",X"0c",X"04",X"08",X"00",X"00",X"00",X"00", 			--  '''
								X"00",X"01",X"02",X"04",X"04",X"04",X"02",X"01", 			--  '('
								X"00",X"08",X"04",X"02",X"02",X"02",X"04",X"08",			--  ')'
								X"00",X"00",X"04",X"15",X"0e",X"15",X"04",X"00", 			--  '*'
								X"00",X"00",X"04",X"04",X"1f",X"04",X"04",X"00", 			--  '+'
								X"00",X"00",X"00",X"00",X"00",X"0c",X"04",X"08", 			--  ','
								X"00",X"00",X"00",X"00",X"1f",X"00",X"00",X"00",			--  '-'
								X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"06", 			--  '.'
								X"00",X"00",X"01",X"02",X"04",X"08",X"10",X"00", 			--  '/'

								X"00",X"0e",X"11",X"13",X"15",X"19",X"11",X"0e",			--  '0'
								X"00",X"04",X"0c",X"04",X"04",X"04",X"04",X"0e",		 	--  '1'
								X"00",X"0e",X"11",X"01",X"02",X"04",X"08",X"1f", 			--  '2'
								X"00",X"1f",X"02",X"04",X"02",X"01",X"11",X"0e",	 		--  '3'
								X"00",X"02",X"06",X"0a",X"12",X"1f",X"02",X"02", 			--  '4'
								X"00",X"1f",X"10",X"1e",X"01",X"01",X"11",X"0e", 			--  '5'
								X"00",X"06",X"08",X"10",X"1e",X"11",X"11",X"0e",	 		--  '6'
								X"00",X"1f",X"01",X"02",X"04",X"08",X"08",X"08",		 	--  '7'
								X"00",X"0e",X"11",X"11",X"0e",X"11",X"11",X"0e",	 		--  '8'
								X"00",X"0e",X"11",X"11",X"0e",X"01",X"02",X"0c",			--  '9'
								X"00",X"00",X"0c",X"0c",X"00",X"0c",X"0c",X"00", 			--  ':'
								X"00",X"00",X"0c",X"0c",X"00",X"0c",X"04",X"08",		 	--  ';'
								X"00",X"02",X"04",X"08",X"10",X"08",X"04",X"02",		 	--  '<'
								X"00",X"00",X"00",X"1f",X"00",X"1f",X"00",X"00",			--  '='
								X"00",X"08",X"04",X"02",X"01",X"02",X"04",X"08", 			--  '>'
								X"00",X"0e",X"11",X"01",X"02",X"04",X"00",X"04", 			--  '?'

								X"00",X"0e",X"11",X"01",X"0d",X"15",X"15",X"0e",	 		--  '@'
								X"00",X"0e",X"11",X"11",X"1f",X"11",X"11",X"11", 			--  'A'
								X"00",X"1e",X"11",X"11",X"1e",X"11",X"11",X"1e", 			--  'B'
								X"00",X"0e",X"11",X"10",X"10",X"10",X"11",X"0e", 			--  'C'
								X"00",X"1c",X"12",X"11",X"11",X"11",X"12",X"1c", 			--  'D'
								X"00",X"1f",X"10",X"10",X"1e",X"10",X"10",X"1f", 			--  'E'
								X"00",X"1f",X"10",X"10",X"1e",X"10",X"10",X"10", 			--  'F'
								X"00",X"0e",X"11",X"10",X"17",X"11",X"11",X"0e", 			--  'G'
								X"00",X"11",X"11",X"11",X"1f",X"11",X"11",X"11", 			--  'H'
								X"00",X"1f",X"04",X"04",X"04",X"04",X"04",X"1f",			--  'I'
								X"00",X"0f",X"02",X"02",X"02",X"02",X"12",X"0c", 			--  'J'
								X"00",X"11",X"12",X"14",X"18",X"14",X"12",X"11", 			--  'K'
								X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"1F", 			--  'L'
								X"00",X"11",X"1B",X"15",X"15",X"11",X"11",X"11",			--  'M'
								X"00",X"11",X"11",X"19",X"15",X"13",X"11",X"11", 			--  'N'
								X"00",X"0e",X"11",X"11",X"11",X"11",X"11",X"0e", 			--  'O'
								X"00",X"1e",X"11",X"11",X"1e",X"10",X"10",X"10", 			--  'P'
								X"00",X"0e",X"11",X"11",X"11",X"15",X"12",X"0d", 			--  'Q'
								X"00",X"1e",X"11",X"11",X"1e",X"14",X"12",X"11", 			--  'R'
								X"00",X"0f",X"10",X"10",X"0e",X"01",X"01",X"1e", 			--  'S'
								X"00",X"1f",X"04",X"04",X"04",X"04",X"04",X"04",		 	--  'T'
								X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"0e", 			--  'U'
								X"00",X"11",X"11",X"11",X"11",X"11",X"0a",X"04",			--  'V'
								X"00",X"11",X"11",X"11",X"11",X"15",X"15",X"0a",			--  'W'
								X"00",X"11",X"11",X"0a",X"04",X"0a",X"11",X"11",	 		--  'X'
								X"00",X"11",X"11",X"11",X"0a",X"04",X"04",X"04",	 		--  'Y'
								X"00",X"1f",X"01",X"02",X"04",X"08",X"10",X"1f",			--  'Z'
								X"00",X"0e",X"08",X"08",X"08",X"08",X"08",X"0e",	 		--  '['
								X"00",X"00",X"10",X"08",X"04",X"02",X"01",X"00",			--  '\'
								X"00",X"0e",X"02",X"02",X"02",X"02",X"02",X"0e",		 	--  ']'
								X"00",X"04",X"0a",X"11",X"00",X"00",X"00",X"00", 			--  '^'
								X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1f",			--  '_'
								X"00",X"08",X"04",X"02",X"00",X"00",X"00",X"00",	 		--  '`'
								
								X"00",X"00",X"00",X"0e",X"01",X"0f",X"11",X"0f",			--  'a'
								X"00",X"10",X"10",X"10",X"1e",X"11",X"11",X"1e", 			--  'b'
								X"00",X"00",X"00",X"0f",X"10",X"10",X"10",X"0f", 			--  'c'
								X"00",X"01",X"01",X"01",X"0f",X"11",X"11",X"0f",	 		--  'd'
								X"00",X"00",X"00",X"0e",X"11",X"1f",X"10",X"0e",		 	--  'e'
								X"00",X"02",X"05",X"04",X"0e",X"04",X"04",X"04", 			--  'f'
								X"00",X"00",X"00",X"0f",X"11",X"0f",X"01",X"1e",		 	--  'g'
								X"00",X"10",X"10",X"10",X"1e",X"11",X"11",X"11", 			--  'h'
								X"00",X"00",X"04",X"00",X"04",X"04",X"04",X"04",			--  'i'
								X"00",X"02",X"00",X"02",X"02",X"02",X"12",X"0c", 			--  'j'
								X"00",X"08",X"08",X"09",X"0a",X"0c",X"0a",X"09",		 	--  'k'
								X"00",X"0c",X"04",X"04",X"04",X"04",X"04",X"0e",		 	--  'l'
								X"00",X"00",X"00",X"1b",X"15",X"15",X"15",X"11",			--  'm'
								X"00",X"00",X"00",X"16",X"19",X"11",X"11",X"11", 			--  'n'
								X"00",X"00",X"00",X"0e",X"11",X"11",X"11",X"0e",	 		--  'o'
								X"00",X"00",X"00",X"1e",X"11",X"1e",X"10",X"10", 			--  'p'
								X"00",X"00",X"00",X"0f",X"11",X"0f",X"01",X"01",		 	--  'q'
								X"00",X"00",X"00",X"16",X"19",X"10",X"10",X"10", 			--  'r'
								X"00",X"00",X"00",X"0f",X"10",X"0e",X"01",X"1e", 			--  's'
								X"00",X"04",X"04",X"1f",X"04",X"04",X"05",X"02",		 	--  't'
								X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"0e", 			--  'u'
								X"00",X"00",X"00",X"11",X"11",X"11",X"0a",X"04",			--  'v'
								X"00",X"00",X"00",X"11",X"11",X"15",X"15",X"0a",			--  'w'
								X"00",X"00",X"00",X"11",X"0a",X"04",X"0a",X"11",	 		--  'x'
								X"00",X"00",X"00",X"11",X"0a",X"04",X"04",X"08",		 	--  'y'
								X"00",X"00",X"00",X"1f",X"02",X"04",X"08",X"1f",			--  'z'
								X"00",X"03",X"04",X"04",X"08",X"04",X"04",X"03",			--  '{'
								X"00",X"04",X"04",X"04",X"00",X"04",X"04",X"04",		 	--  '|'
								X"00",X"18",X"04",X"04",X"03",X"04",X"04",X"18",	 		--  ''
								X"00",X"00",X"08",X"15",X"02",X"00",X"00",X"00",			--  '~'
								others => X"00"
						);
Begin
	process(Address)
		variable	index : integer range 0 to 1023 ;	
	begin
		index := to_integer(unsigned(Address)) ;
		DataOut <= MyRom(index);
	end process ;
END ;

