library verilog;
use verilog.vl_types.all;
entity MC68K_vlg_vec_tst is
end MC68K_vlg_vec_tst;
