library verilog;
use verilog.vl_types.all;
entity MC68K_vlg_check_tst is
    port(
        Address_OUT     : in     vl_logic_vector(31 downto 0);
        AddressBus      : in     vl_logic_vector(31 downto 0);
        AS_L            : in     vl_logic;
        AS_OUT_L        : in     vl_logic;
        BG_L            : in     vl_logic;
        BGACK_L         : in     vl_logic;
        BlueOut         : in     vl_logic_vector(9 downto 0);
        BR_L            : in     vl_logic;
        CPU_RW          : in     vl_logic;
        CPUClock        : in     vl_logic;
        DataBusIn       : in     vl_logic_vector(15 downto 0);
        DataBusOut      : in     vl_logic_vector(15 downto 0);
        DMA_DataOut     : in     vl_logic_vector(15 downto 0);
        DramDtack_L     : in     vl_logic;
        DramSelect_H    : in     vl_logic;
        Dtack_L         : in     vl_logic;
        FlashAddress    : in     vl_logic_vector(21 downto 0);
        FlashCE_L       : in     vl_logic;
        FlashData       : in     vl_logic_vector(7 downto 0);
        FlashOE_L       : in     vl_logic;
        FlashReset_L    : in     vl_logic;
        FlashWE_L       : in     vl_logic;
        GreenLEDS       : in     vl_logic_vector(7 downto 0);
        GreenOut        : in     vl_logic_vector(9 downto 0);
        HexDisplay0     : in     vl_logic_vector(6 downto 0);
        HexDisplay1     : in     vl_logic_vector(6 downto 0);
        HexDisplay2     : in     vl_logic_vector(6 downto 0);
        HexDisplay3     : in     vl_logic_vector(6 downto 0);
        HexDisplay4     : in     vl_logic_vector(6 downto 0);
        HexDisplay5     : in     vl_logic_vector(6 downto 0);
        HexDisplay6     : in     vl_logic_vector(6 downto 0);
        HexDisplay7     : in     vl_logic_vector(6 downto 0);
        horiz_sync_out  : in     vl_logic;
        LCD_BLON_DE2    : in     vl_logic;
        LCD_Contrast_DE1: in     vl_logic;
        LCD_E           : in     vl_logic;
        LCD_ON_DE2      : in     vl_logic;
        LCD_RS          : in     vl_logic;
        LCD_RW          : in     vl_logic;
        LCDDataOut      : in     vl_logic_vector(7 downto 0);
        LDS_L           : in     vl_logic;
        LDS_OUT_L       : in     vl_logic;
        OnChipRamSelect_H: in     vl_logic;
        OutPortE        : in     vl_logic_vector(7 downto 0);
        RedLEDSA        : in     vl_logic_vector(7 downto 0);
        RedLEDSB        : in     vl_logic_vector(7 downto 0);
        RedLEDSC        : in     vl_logic_vector(7 downto 0);
        RedOut          : in     vl_logic_vector(9 downto 0);
        ResetOut        : in     vl_logic;
        RomSelect_H     : in     vl_logic;
        RS232_TxData    : in     vl_logic;
        RW_OUT          : in     vl_logic;
        sdram_a         : in     vl_logic_vector(11 downto 0);
        sdram_ba        : in     vl_logic_vector(1 downto 0);
        sdram_cas_n     : in     vl_logic;
        sdram_cke       : in     vl_logic;
        sdram_clock     : in     vl_logic;
        sdram_cs_n      : in     vl_logic;
        sdram_dq        : in     vl_logic_vector(15 downto 0);
        sdram_dqm       : in     vl_logic_vector(1 downto 0);
        sdram_ras_n     : in     vl_logic;
        sdram_we_n      : in     vl_logic;
        SRam_CE_L       : in     vl_logic;
        SRam_Data       : in     vl_logic_vector(15 downto 0);
        SRam_LB_L       : in     vl_logic;
        SRam_OE_L       : in     vl_logic;
        SRam_UB_L       : in     vl_logic;
        SRam_WE_L       : in     vl_logic;
        SRamAddress     : in     vl_logic_vector(17 downto 0);
        SRamSelect_H    : in     vl_logic;
        UDS_L           : in     vl_logic;
        UDS_OUT_L       : in     vl_logic;
        vert_sync_out   : in     vl_logic;
        VideoDAC_Blank_L: in     vl_logic;
        VideoDac_Clock  : in     vl_logic;
        VideoDac_Sync_L : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MC68K_vlg_check_tst;
